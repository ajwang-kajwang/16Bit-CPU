library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity RAM is
  port (
    clk  : in std_logic;
    addr : in std_logic_vector(15 downto 0); -- Changed address width to 8 bits
    data : inout std_logic_vector(15 downto 0);
    we   : in std_logic -- Write enable
  );
end entity;

architecture behavioral of RAM is
  type ram_type is array (0 to 255) of std_logic_vector(15 downto 0);
  signal ram      : ram_type := (others => (others => '0'));
  signal data_out : std_logic_vector(15 downto 0);

begin
  process (clk)
  begin
    if rising_edge(clk) and addr(15 downto 12) = "1000" then
      if we = '1' then
        ram(to_integer(unsigned(addr(7 downto 0)))) <= data;
      else
        data_out <= ram(to_integer(unsigned(addr(7 downto 0))));
      end if;
    end if;
  end process;

  data <= data_out when (we = '0'and addr(15 downto 12) = "1000") else
    (others => 'Z');

end behavioral;